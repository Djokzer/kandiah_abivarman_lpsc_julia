library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity gen_complex is
    port (
        clk   : in std_logic;
        reset : in std_logic
    );
end entity gen_complex;

architecture rtl of gen_complex is

begin

    

end architecture;