library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity julia_compute is
    port (
        clk   : in std_logic;
        reset : in std_logic
        
    );
end entity julia_compute;

architecture rtl of julia_compute is

begin

    

end architecture;